`include ../rtl/include/cv32e40p_pkg.sv

module cv32e40p_alu
 import cv32e40p_pkg::*;
(
    input logic               clk,
    input logic               rst_n,
    input logic               enable_i,
    input alu_opcode_e        operator_i,
    input logic        [31:0] operand_a_i,
    input logic        [31:0] operand_b_i,
	);

endmodule
