package tb_pkg;
	import uvm_pkg::*;

//`include "test_cfg.svh"
//`include "alu_package.svh"
`include "alu_transaction.svh"
`include "alu_sequence.svh"
`include "alu_driver.svh"
`include "alu_seqr.svh"
`include "alu_agent.svh"
//`include "alu_coverage.svh"
`include "alu_env.svh"
`include "alu_test.svh";

endpackage
